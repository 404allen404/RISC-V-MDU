`ifndef MDU_DEFINE
`define MDU_DEFINE 1

`define MD_ALU_ADD 2'b00
`define MD_ALU_SUB 2'b01
`define MD_ALU_NOP 2'b10

`endif